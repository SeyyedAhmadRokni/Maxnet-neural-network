module MUX2(input sel , input[31:0] , a , b , output[31:0] out);
    
endmodule