module  TestBench();
    reg clk=0 ,start=0 ,rst=0;
    reg [31:0] eps=32'b10111110010011001100110011001101 ,
    a1 = 32'b01000010111111010110011001100110,
    a2 = 32'b11000000101000000000000000000000,
    a3 = 32'b00000000000000000000000000000000,
    a4 = 32'b10111110010011001100110011001101;
    always #5 clk = ~clk;
    wire finish;
    wire [31 : 0] out;
    // reg[31:0] x1 = 32'b01000010111111010110011001100110,x2 = 32'b11000000101000000000000000000000 //12..  -5
    // ,x3 = 32'b00000000000000000000000000000000,x4 = 32'b01000010101010110110000101001000  // 0   85...
    // , e = 32'b10111110010011001100110011001101; // -0.2
    Maxnet_model mxn( start , clk ,eps , a1 , a2 , a3 , a4 ,  finish , out);
    initial begin
        #12 start=1;
        #10 start=0;

        #2000 
        $stop;
    end

endmodule