module Mul_test();
    reg [31:0] a, b;
    reg clk = 1'b0;
    wire [31:0] out;
    Mul ml(a, b, out);
    always begin
        #5;
        clk = ~clk;
    end

    initial begin
        a = 32'b00111111110000010100011110101110; //1.51
        b = 32'b01000000001101010001111010111000; //2.83
        #40;
        b = 32'b01000000011010011001100110011010; //3.65
        #40;
        a = 32'b00000000000000000000000000000000; //0
        b = 32'b00000000000000000000000000000000; //0
        #40;

        $stop;

    end


endmodule